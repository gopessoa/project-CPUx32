module cpu(
    input wire clk,
    input wire reset
);

endmodule